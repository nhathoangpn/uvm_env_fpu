//==================================================================================================
// Owner:    Hoang Pham
// Filename: fpu_test_pkg
// History:  2019.06.21 Create new version
//==================================================================================================

package fpu_test_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	import fpu_env_pkg::*;
	import fpu_agent_pkg::*;

	`include "fpu_test_base.sv"

	`include "fpu_test_sample_00.sv"
	`include "fpu_test_sample_01.sv"
	`include "fpu_test_sample_02.sv"
	`include "fpu_test_sample_03.sv"
	`include "fpu_test_sample_04.sv"
	`include "fpu_test_sample_05.sv"

	// list all test scenarios here
	`include "fpu_error_test_arth.sv"
	`include "fpu_error_test_cmpcvt.sv"
	`include "fpu_error_test_dis_arth.sv"
	`include "fpu_error_test_dis_cmpcvt.sv"
	`include "fpu_error_test_dis_explog.sv"
	`include "fpu_error_test_dis_sm.sv"
	`include "fpu_error_test_reserved_pipeline.sv"
	`include "fpu_error_test_sm.sv"
	`include "fpu_para_test_en_all_dis_explog.sv"
	`include "fpu_para_test_en_all_en_explog.sv"
	`include "fpu_para_test_en_arth_cmpcvt.sv"
	`include "fpu_para_test_en_arth_sm_dis_explog.sv"
	`include "fpu_para_test_en_arth_sm_en_explog.sv"
	`include "fpu_para_test_en_arth.sv"
	`include "fpu_para_test_en_cmpcvt_sm_dis_explog.sv"
	`include "fpu_para_test_en_cmpcvt_sm_en_explog.sv"
	`include "fpu_para_test_en_cmpcvt.sv"
	`include "fpu_para_test_en_sm_dis_explog.sv"
	`include "fpu_para_test_en_sm_en_explog.sv"
	`include "fpu_test_add.sv"
	`include "fpu_test_add_u.sv"
	`include "fpu_test_arth_sm_compcvt_invld.sv"
	`include "fpu_test_arth_sm_compcvt_vld.sv"
	`include "fpu_test_conflict_stall_reset.sv"
	`include "fpu_test_div_s.sv"
	`include "fpu_test_div_u.sv"
	`include "fpu_test_fadd.sv"
	`include "fpu_test_fcvt_s_w.sv"
	`include "fpu_test_fcvt_s_wu.sv"
	`include "fpu_test_fcvt_w_s.sv"
	`include "fpu_test_fcvt_wu_s.sv"
	`include "fpu_test_fdiv.sv"
	`include "fpu_test_feq.sv"
	`include "fpu_test_fexp.sv"
	`include "fpu_test_fle.sv"
	`include "fpu_test_flog.sv"
	`include "fpu_test_flt.sv"
	`include "fpu_test_fmadd.sv"
	`include "fpu_test_fmax.sv"
	`include "fpu_test_fmin.sv"
	`include "fpu_test_fmnadd.sv"
	`include "fpu_test_fmnsub.sv"
	`include "fpu_test_fmsub.sv"
	`include "fpu_test_fmul.sv"
	`include "fpu_test_fne.sv"
	`include "fpu_test_fsqrt.sv"
	`include "fpu_test_fsub.sv"
	`include "fpu_test_input_flush_fadd.sv"
	`include "fpu_test_input_flush_fcvt_w_s.sv"
	`include "fpu_test_input_flush_fcvt_wu_s.sv"
	`include "fpu_test_input_flush_fdiv.sv"
	`include "fpu_test_input_flush_feq.sv"
	`include "fpu_test_input_flush_fexp.sv"
	`include "fpu_test_input_flush_fle.sv"
	`include "fpu_test_input_flush_flog.sv"
	`include "fpu_test_input_flush_flt.sv"
	`include "fpu_test_input_flush_fmadd.sv"
	`include "fpu_test_input_flush_fmax.sv"
	`include "fpu_test_input_flush_fmin.sv"
	`include "fpu_test_input_flush_fmnadd.sv"
	`include "fpu_test_input_flush_fmnsub.sv"
	`include "fpu_test_input_flush_fmsub.sv"
	`include "fpu_test_input_flush_fmul.sv"
	`include "fpu_test_input_flush_fne.sv"
	`include "fpu_test_input_flush_fsqrt.sv"
	`include "fpu_test_input_flush_fsub.sv"
	`include "fpu_test_madd.sv"
	`include "fpu_test_mnadd.sv"
	`include "fpu_test_mnsub.sv"
	`include "fpu_test_msub.sv"
	`include "fpu_test_mulh_su.sv"
	`include "fpu_test_mulh.sv"
	`include "fpu_test_mulh_u.sv"
	`include "fpu_test_mul_su.sv"
	`include "fpu_test_mul.sv"
	`include "fpu_test_mul_u.sv"
	`include "fpu_test_nonpipeline_sm_invld.sv"
	`include "fpu_test_nonpipeline_sm_vld.sv"
	`include "fpu_test_output_flush_fadd.sv"
	`include "fpu_test_output_flush_fdiv.sv"
	`include "fpu_test_output_flush_fexp.sv"
	`include "fpu_test_output_flush_flog.sv"
	`include "fpu_test_output_flush_fmadd.sv"
	`include "fpu_test_output_flush_fmnadd.sv"
	`include "fpu_test_output_flush_fmnsub.sv"
	`include "fpu_test_output_flush_fmsub.sv"
	`include "fpu_test_output_flush_fmul.sv"
	`include "fpu_test_output_flush_fsqrt.sv"
	`include "fpu_test_output_flush_fsub.sv"
	`include "fpu_test_pipeline_arth_cmpcvt.sv"
	`include "fpu_test_pipeline_arth.sv"
	`include "fpu_test_pipeline_cmpcvt.sv"
	`include "fpu_test_rem_s.sv"
	`include "fpu_test_rem_u.sv"
	`include "fpu_test_rst_arth.sv"
	`include "fpu_test_rst_cmpcvt.sv"
	`include "fpu_test_rst_init_error_o.sv"
	`include "fpu_test_rst_init.sv"
	`include "fpu_test_rst_sm.sv"
	`include "fpu_test_stall_arth.sv"
	`include "fpu_test_stall_cmpcvt.sv"
	`include "fpu_test_stall_rand.sv"
	`include "fpu_test_stall_sm.sv"
	`include "fpu_test_sub.sv"
	`include "fpu_test_sub_u.sv"

	`include "fpu_test_fsqrt_all_man.sv"
	`include "fpu_test_flog_all_man.sv"
	`include "fpu_test_fexp_all_man.sv"

	`include "fpu_test_reserved_rm.sv"

	// list all direct debug test scenarios here
	`include "debug_test/fpu_test_fadd_db_3457_01.sv"
	`include "debug_test/fpu_test_fadd_db_3457_02.sv"
	`include "debug_test/fpu_test_fadd_db_3457_03.sv"
	`include "debug_test/fpu_test_fadd_db_3458_01.sv"
	`include "debug_test/fpu_test_fadd_db_3504_01.sv"
	`include "debug_test/fpu_test_fdiv_db_3505_01_inf_p.sv"
	`include "debug_test/fpu_test_fdiv_db_3505_02_inf_m.sv"
	`include "debug_test/fpu_test_fdiv_db_3505_03_zero_p.sv"
	`include "debug_test/fpu_test_fdiv_db_3505_04_zero_m.sv"
	`include "debug_test/fpu_test_fdiv_db_3505_05_cNAN.sv"
	`include "debug_test/fpu_test_fdiv_db_3505_06_A_zero.sv"
	`include "debug_test/fpu_test_fdiv_db_3505_07_A_sn.sv"
	`include "debug_test/fpu_test_fdiv_db_3505_08_B_sn.sv"
	`include "debug_test/fpu_test_fdiv_db_3505.sv"
	`include "debug_test/fpu_test_fexp_db_3525.sv"
	`include "debug_test/fpu_test_flog_db_3485_01.sv"
	`include "debug_test/fpu_test_flog_db_3485_02.sv"
	`include "debug_test/fpu_test_flog_db_3485_03.sv"
	`include "debug_test/fpu_test_fmadd_db_01.sv"
	`include "debug_test/fpu_test_fmadd_db_spec_3495_01.sv"
	`include "debug_test/fpu_test_fmul_db_3460_01.sv"
	`include "debug_test/fpu_test_fmul_db_3506.sv"
	`include "debug_test/fpu_test_fmul_db_3508.sv"
	`include "debug_test/fpu_test_fsqrt_all_man_db_3514_01.sv"
	`include "debug_test/fpu_test_mul_db_3517.sv"
	`include "debug_test/fpu_test_mulh_db_3519.sv"
	`include "debug_test/fpu_test_mulh_u_db_3520.sv"
	`include "debug_test/fpu_test_sub_db_3516.sv"
	`include "debug_test/fpu_test_fsqrt_db_3489_01_case1.sv"
	`include "debug_test/fpu_test_add_db_3486.sv"
	`include "debug_test/fpu_test_div_db_3487.sv"
	`include "debug_test/fpu_test_div_u_db_3488.sv"
	`include "debug_test/fpu_test_madd_db_3490.sv"
	`include "debug_test/fpu_test_mnadd_db_3490.sv"
	`include "debug_test/fpu_test_msub_db_3490.sv"
	`include "debug_test/fpu_test_mnsub_db_3490.sv"
	`include "debug_test/fpu_test_mul_db_3499.sv"
	`include "debug_test/fpu_test_mulh_db_3499.sv"
	`include "debug_test/fpu_test_flog_db_3500.sv"
	`include "debug_test/fpu_test_rem_db_3529.sv"
	`include "debug_test/fpu_test_rem_u_db_3529.sv"
	`include "debug_test/fpu_test_flog_man_a_fix_1_0000xxxx.sv"
	`include "debug_test/fpu_test_flog_man_a_fix_2_0000xxxx.sv"
	`include "debug_test/fpu_test_flog_man_a_fix_7E_7FFFxx.sv"
	`include "debug_test/fpu_test_flog_man_a_fix_7E_7Fxxxx.sv"
	`include "debug_test/fpu_test_flog_man_a_fix_7E_xxxxxx.sv"
    `include "fpu_test_fexp_negative_int.sv"
    `include "fpu_test_fexp_positive_int.sv"
    `include "fpu_test_fexp_sub_normal.sv"
    `include "fpu_test_fexp_negative_126.sv"
    `include "fpu_test_fexp_negative_127.sv"
    `include "fpu_test_fexp_zero.sv"
    `include "fpu_test_flog_1_0.sv"
    `include "fpu_test_flog_sub_normal.sv"
    `include "debug_test/fpu_test_flog_1_5_to_2_0.sv"
    `include "debug_test/fpu_test_flog_0_5_to_1_0.sv"
    `include "debug_test/fpu_test_flog_1_0_to_1_5.sv"


	// list all ccov improving scenarios here
	`include "fpu_test_div_dz_cov_improve.sv"
	`include "fpu_test_div_u_dz_cov_improve.sv"
	`include "fpu_test_rem_dz_cov_improve.sv"
	`include "fpu_test_rem_u_dz_cov_improve.sv"
	`include "fpu_test_fmadd_unf_1_cov_improve.sv"
	`include "fpu_test_fmadd_unf_2_cov_improve.sv"
	`include "fpu_test_flog_man_a_zero_cov_improve.sv"
	`include "fpu_test_cnv_cov_improve.sv"
	`include "fpu_test_packed_cov_improve.sv"
	`include "fpu_test_fsqrt_SRT_cov_improve.sv"
	`include "fpu_test_fexp_norm_cov_improve.sv"
	`include "fpu_test_flog_cnt_pointer_cov_improve.v"
	`include "fpu_test_none_calc_cov_improve.v"
	`include "fpu_test_fcov_uf_of_fmadd.sv"
	`include "fpu_test_fcov_fexp_grs_010_100_110.sv"
	`include "fpu_test_arith_ccov_improve.sv"
	`include "fpu_test_fcov_flog_lzc.sv"

	// list all fcov improving scenarios here
	`include "fpu_test_fcov_rst_during_calc.sv"
	`include "fpu_test_fcov_round_w_output_flushing.sv"
	`include "fpu_test_fcov_stall_reset_type1.sv"
	`include "fpu_test_fcov_stall_reset_type2.sv"
	`include "fpu_test_fcov_cs_op_operand.sv"
	`include "fpu_test_fcov_fcvt_w_wu_s_out_of_range.sv"
	`include "fpu_test_fcov_nx_0.sv"
	`include "fpu_test_fcov_cg_FPU_Flags_Coverage.sv"
	`include "fpu_test_fcov_cg_Result_format_Arith_fmxxx.sv"

	//For GRS fcov
	`include "fpu_test_fcov_fmul_grs_xx0.sv"

endpackage
