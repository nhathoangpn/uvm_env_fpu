//==================================================================================================
// Owner:    Thinh.Le
// Filename: fpu_test_fcov_fmul_grs_xx0
// History:  2019.10.24 Create new version
//==================================================================================================

class fpu_test_fcov_fmul_grs_xx0 extends fpu_test_base;
	`uvm_component_utils(fpu_test_fcov_fmul_grs_xx0)

	`include "../fpu_top/fpu_def.svh"

	fpu_seq_base seq_srandom;
	fpu_seq_base seq_final;

	function new(string name, uvm_component parent);
		super.new(name, parent);
	endfunction

	task run_phase(uvm_phase phase);
		phase.phase_done.set_drain_time(this, 110);
		phase.raise_objection(this, {get_name, "run_phase starts"});
		`uvm_info(get_name(), "run_phase starts", UVM_FULL)

		m_fpu_agent_cfg.fpu_vif.rst_gen_direct(1, 10);

		seq_srandom = fpu_seq_base::type_id::create("seq_srandom");
		seq_final   = fpu_seq_base::type_id::create("seq_final");

		for (int i = 0; i < 1000; i++) begin
			for (int j = 0; j < 5; j++) begin
				if (!seq_srandom.randomize() with
					{sub_num_seq_item == 1;
					 sqb_valid_i == 1;
					 sqb_op_i == `FMUL;
					 sqb_operand_b_i[20:0] == 21'h0;
					 sqb_rm_i == j;
					 sqb_fn_i == 0;
					 sqb_user_i inside{[8'h00:8'hFF]};
					 sqb_num_wait_clk == 1;
					 sqb_test_final == 0;
					 sqb_handshake_i == 0;
					})
				`uvm_error("RANDOM SEQUENCE", "randomization failure for sequence")

				seq_srandom.start(m_fpu_env.m_fpu_agent.m_fpu_sqr);
			end
		end

		if (!seq_final.randomize() with
			{sub_num_seq_item == 1;
			 sqb_num_wait_clk == 1;
			 sqb_test_final   == 1;})
		`uvm_error("FINAL SEQUENCE", "randomization failure for sequence")

		seq_final.start(m_fpu_env.m_fpu_agent.m_fpu_sqr);

		phase.drop_objection(this, {get_name, "run_phase finishes"});
		`uvm_info(get_name(), "run_phase finishes", UVM_FULL)
	endtask
endclass
