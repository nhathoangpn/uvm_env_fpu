//==================================================================================================
// Owner:    Hoang Pham
// Filename: fpu_env_pkg
// History:  2019.06.21 Create new version
//==================================================================================================

package fpu_env_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	import fpu_agent_pkg::*;

	`include "fpu_env_cfg.sv"
	`include "fpu_scb.sv"
	`include "fpu_fcov.sv"
	`include "fpu_env.sv"
endpackage
