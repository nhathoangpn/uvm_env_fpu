//==================================================================================================
// Owner:    Thinh Le
// Filename: for fcov
// History:  2019.06.21 Create new version
//==================================================================================================

class fpu_test_fcov_fcvt_w_wu_s_out_of_range extends fpu_test_base;
	`uvm_component_utils(fpu_test_fcov_fcvt_w_wu_s_out_of_range)

	`include "../fpu_top/fpu_def.svh"

	fpu_seq_base seq_srandom;
	fpu_seq_base seq_sdirect;
	fpu_seq_base seq_final;

	function new(string name, uvm_component parent);
		super.new(name, parent);
	endfunction

	task run_phase(uvm_phase phase);
		phase.phase_done.set_drain_time(this, 110);
		phase.raise_objection(this, {get_name, "run_phase starts"});
		`uvm_info(get_name(), "run_phase starts", UVM_FULL)

		m_fpu_agent_cfg.fpu_vif.rst_gen_direct(1, 10);

		seq_srandom = fpu_seq_base::type_id::create("seq_srandom");
		seq_sdirect = fpu_seq_base::type_id::create("seq_sdirect");
		seq_final   = fpu_seq_base::type_id::create("seq_final");

		for (int i = 0; i < 100; i++) begin
			for (int j = 0; j < 5; j++) begin
				if (!seq_srandom.randomize() with
					{sub_num_seq_item == 1;
					 sqb_valid_i == 1;
					 sqb_op_i inside {`FCVT_W_S, `FCVT_WU_S};
					 sqb_operand_a_i inside {32'h4EFF_FFFF, 32'h4F00_0000, 32'hCEFF_FFFF,  32'hCF00_0000, 32'hCF00_0001, 32'h4F7F_FFFF, 32'h4F80_0000};
					 sqb_rm_i == j;
					 sqb_fn_i == 0;
					 sqb_user_i inside{[8'h00:8'hFF]};
					 sqb_num_wait_clk == 1;
					 sqb_test_final == 0;
					 sqb_handshake_i == 1;})
				`uvm_error("RANDOM SEQUENCE", "randomization failure for sequence")
	
				seq_srandom.start(m_fpu_env.m_fpu_agent.m_fpu_sqr);
			end
		end

		if (!seq_final.randomize() with
			{sub_num_seq_item == 1;
			 sqb_num_wait_clk == 1;
			 sqb_test_final   == 1;})
		`uvm_error("RANDOM SEQUENCE", "randomization failure for sequence")

		seq_final.start(m_fpu_env.m_fpu_agent.m_fpu_sqr);

		phase.drop_objection(this, {get_name, "run_phase finishes"});
		`uvm_info(get_name(), "run_phase finishes", UVM_FULL)
	endtask
endclass
